* C:\SPB_Data\eSim-Workspace\anand_seq\anand_seq.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10-Mar-22 7:02:30 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ Net-_U4-Pad4_ anand_seq		
U5  Net-_U1-Pad~_ Net-_U2-Pad~_ Net-_U3-Pad~_ Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ adc_bridge_3		
U6  Net-_U4-Pad4_ Net-_R1-Pad1_ adc_bridge_1		
v1  Net-_U1-Pad~_ GND pulse		
v2  Net-_U2-Pad~_ GND pulse		
v3  Net-_U3-Pad~_ GND pulse		
U1  Net-_U1-Pad~_ plot_v1		
U2  Net-_U2-Pad~_ plot_v1		
U3  Net-_U3-Pad~_ plot_v1		
U7  out plot_v1		
R1  Net-_R1-Pad1_ out 1k		
C1  out GND 1u		

.end
